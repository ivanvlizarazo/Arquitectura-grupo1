library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity InstructionMemory is
port (
		rst: in std_logic;
      Addr : in std_logic_vector(31 downto 0);
      Instruction : out std_logic_vector(31 downto 0));
end InstructionMemory;

architecture syn of InstructionMemory is
    type rom_type is array (0 to 63) of std_logic_vector (31 downto 0);                 
    signal ROM : rom_type:= ("00000000000000000000000000000000",
										"10100000000100000010000000000110",
"10100010000100000010000000000100",
"10100100000100000010000000000000",
"10100110000100000010000000000001",
"10000000101001000110000000000000",
"00000010100000000000000000001101",
"00000000000000000000000000000000",
"01000000000000000000000000000100",
"00000000000000000000000000000000",
"00010000100000000000000000001010",
"00000000000000000000000000000000",
"10101000000001001000000000010000",
"10100100000100000000000000010100",
"10000000101001001100000000010001",
"10101010000001001110000000000001",
"00001100101111111111111111111100",
"10100110000100000000000000010101",
"10000001110000111110000000000010",
"10010000000100000000000000010010",
"10010000000100000010000000000000",
"00000000000000000000000000000000",
									  others => "00000000000000000000000000000000"); 
begin
    process (rst, Addr)
    begin
		if (rst = '1') then
			Instruction <= "00000000000000000000000000000000";
      else 
			Instruction <= ROM(conv_integer(Addr));
		end if;
    end process;

end syn;

